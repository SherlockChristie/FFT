
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);




    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = 1'b0;
    assign module_intf_1.ap_ready = 1'b0;
    assign module_intf_1.ap_done = 1'b0;
    assign module_intf_1.ap_continue = 1'b0;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;

    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_ST_fsm_state1;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_ST_fsm_state1;
    assign upc_loop_intf_1.quit_state = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_ST_fsm_state1;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_1.quit_block = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_1.iter_start_enable = 1'b1;
    assign upc_loop_intf_1.iter_end_enable = 1'b1;
    assign upc_loop_intf_1.quit_enable = 1'b1;
    assign upc_loop_intf_1.loop_start = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_fft32.grp_fft32_Pipeline_input_loop_fu_332.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_2.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_2.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_402.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_3.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_3.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_410.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(1) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_4.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_4.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_418.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(1) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_5.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_5.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_426.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_6.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_6.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_434.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b1;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_7.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_7.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_447.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_8.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_8.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_455.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_9.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_9.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_463.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_10.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_10.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_471.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_11.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_11.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_479.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;
    upc_loop_intf#(1) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_12.quit_enable = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_12.loop_start = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_fft32.grp_generic_sincos_16_4_s_fu_487.grp_generic_sincos_16_4_Pipeline_VITIS_LOOP_87_1_fu_73.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(1) upc_loop_monitor_12;
    upc_loop_intf#(1) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.quit_state = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.quit_enable = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.loop_start = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_fft32.grp_fft32_Pipeline_output_loop_fu_495.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b1;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(1) upc_loop_monitor_13;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);




    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
